module frequency_divider_cpu(input logic clk, reset, output logic clk_out);	

	logic [24:0] counter;

	always_ff @(posedge clk, posedge reset)
		begin
			if(reset)
				begin
					counter <= 25'd0;
					clk_out <= 1'b0;
				end
			else if(counter == 25'd12500000)
				begin
					counter <= 25'd0;
					clk_out <= ~clk_out;
				end
			else
				begin
					counter <= counter + 1'b1;
				end
		end

endmodule

