module Sprite(input logic [9:0] posX, posY, pixelX, pixelY, output logic [23:0] RGB, output logic isActive);

	logic [1:0] codedColor;
	logic hActive, vActive;

	logic [1:0] sprite [0:31][0:31] =
		'{
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}
		 };

	 assign codedColor = sprite[pixelX - posX][pixelY - posY];
	 
	 decoRGB deco(codedColor, RGB);
	 
	 assign hActive = ((pixelX == posX) || (pixelX < (posX + 32)));
	 assign vActive = ((pixelY == posY) || (pixelY < (posY + 32)));
	
	 assign isActive = hActive & vActive;
	 

endmodule 