module Sprite(input logic [9:0] posX, posY, pixelX, pixelY, input logic [1:0] selec, output logic [23:0] RGB, output logic isActive);

	logic [1:0] codedColorSprite;
	logic [1:0] codedColorSprite1;
	logic [1:0] codedColorSprite2;
	logic [1:0] codedColorSprite3;
	
	logic [1:0] codedColor;
	
	logic hActive, vActive;

	logic [1:0] sprite [0:31][0:31] =
		'{
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
		'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}
		 };
		 
	 logic [1:0] sprite1 [0:31][0:31] =
	'{
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}
	};
		 
	 logic [1:0] sprite2 [0:31][0:31] =
	'{
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}
	};
		 
	 logic [1:0] sprite3 [0:31][0:31] =
	'{
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b10, 2'b10, 2'b11, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}, 
	'{2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01}
	};
	
	 assign codedColorSprite = sprite[pixelX - posX][pixelY - posY];
	 assign codedColorSprite1 = sprite1[pixelX - posX][pixelY - posY];
	 assign codedColorSprite2 = sprite2[pixelX - posX][pixelY - posY];
	 assign codedColorSprite3 = sprite3[pixelX - posX][pixelY - posY];
	 
	 mux_4_x_1 #(2) mux0(codedColorSprite, codedColorSprite1, codedColorSprite2, codedColorSprite3, selec, codedColor); 
	 
	 decoRGB deco(codedColor, RGB);
	 
	 assign hActive = ((pixelX > posX) & (pixelX < (posX + 32)));
	 assign vActive = ((pixelY > posY) & (pixelY < (posY + 25)));
	
	 assign isActive = hActive & vActive;
	 

endmodule 