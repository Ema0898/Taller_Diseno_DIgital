module alu_deco(input logic [3:0] cmd, output logic [3:0] alu_control);

	always_comb
		case(cmd)		
			4'b0000: 
				alu_control = 4'b1000;				
			4'b0001:
				alu_control = 4'b1010;	
			4'b0010:
				alu_control = 4'b0001;
			4'b0100:
				alu_control = 4'b0000;
			4'b1010:
				alu_control = 4'b0001;
			4'b1011:
				alu_control = 4'b0000;
			4'b1100:
				alu_control = 4'b1001;
			4'b1111:
				alu_control = 4'b1011;
		default:
				alu_control = 4'b0000;			
		endcase

endmodule 