module processor(input logic clk,
					  input logic rst,
					  input logic [31:0] instruction, read_data,
					  output logic [31:0] pc, direction, write_data,
					  output logic mem_write);
					  

endmodule 