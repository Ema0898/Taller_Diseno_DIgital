module reg_file_deco(input logic [3:0] x, output logic [15:0] y);

endmodule 