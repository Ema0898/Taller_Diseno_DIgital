module Enemy(input logic [9:0] posX, posY, pixelX, pixelY, output logic [23:0] RGB, output logic isActive);

  logic [2:0] codedColorSprite;	
	
  logic hActive, vActive;

  logic [2:0] sprite [0:31][0:31] =
  '{
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}
};
	
	
	
  assign codedColorSprite = sprite[pixelX - posX][pixelY - posY];
	 	 
  decoRGBEnemy deco(codedColorSprite, RGB);
	 
  assign hActive = ((pixelX > posX) & (pixelX < (posX + 32)));
  assign vActive = ((pixelY > posY) & (pixelY < (posY + 32)));
	
  assign isActive = hActive & vActive; 



endmodule 